magic
tech sky130A
magscale 1 2
timestamp 1713341356
<< nwell >>
rect 3796 1524 6132 1720
rect 3800 -432 6132 1524
<< mvndiff >>
rect 5654 -606 5666 -562
<< mvpsubdiff >>
rect 3210 -656 3252 -632
rect 3210 -722 3252 -698
rect 3210 -913 3252 -889
rect 3210 -979 3252 -955
rect 3210 -1170 3252 -1146
rect 3210 -1236 3252 -1212
rect 3210 -1428 3252 -1404
rect 3210 -1494 3252 -1470
<< mvnsubdiff >>
rect 4198 1630 4240 1654
rect 4198 1564 4240 1588
rect 4574 1630 4616 1654
rect 4574 1564 4616 1588
rect 4950 1630 4992 1654
rect 4950 1564 4992 1588
rect 5326 1630 5368 1654
rect 5326 1564 5368 1588
rect 5702 1630 5744 1654
rect 5702 1564 5744 1588
<< mvpsubdiffcont >>
rect 3210 -698 3252 -656
rect 3210 -955 3252 -913
rect 3210 -1212 3252 -1170
rect 3210 -1470 3252 -1428
<< mvnsubdiffcont >>
rect 4198 1588 4240 1630
rect 4574 1588 4616 1630
rect 4950 1588 4992 1630
rect 5326 1588 5368 1630
rect 5702 1588 5744 1630
<< locali >>
rect 4198 1630 4240 1646
rect 4198 1572 4240 1588
rect 4574 1630 4616 1646
rect 4574 1572 4616 1588
rect 4950 1630 4992 1646
rect 4950 1572 4992 1588
rect 5326 1630 5368 1646
rect 5326 1572 5368 1588
rect 5702 1630 5744 1646
rect 5702 1572 5744 1588
rect 3210 -656 3252 -640
rect 3210 -714 3252 -698
rect 3210 -913 3252 -897
rect 3210 -971 3252 -955
rect 3210 -1170 3252 -1154
rect 3210 -1228 3252 -1212
rect 3210 -1428 3252 -1412
rect 3210 -1486 3252 -1470
<< viali >>
rect 4198 1588 4240 1630
rect 4574 1588 4616 1630
rect 4950 1588 4992 1630
rect 5326 1588 5368 1630
rect 5702 1588 5744 1630
rect 3210 -698 3252 -656
rect 3210 -955 3252 -913
rect 3210 -1212 3252 -1170
rect 3210 -1470 3252 -1428
<< metal1 >>
rect 3204 1272 3442 1704
rect 3536 1272 3774 1704
rect 4186 1653 5756 1691
rect 4186 1636 4252 1653
rect 3874 1458 4046 1590
rect 4186 1584 4193 1636
rect 4245 1584 4252 1636
rect 4562 1630 4628 1653
rect 4562 1588 4574 1630
rect 4616 1588 4628 1630
rect 4938 1630 5004 1653
rect 4682 1603 4874 1610
rect 4682 1590 4694 1603
rect 4186 1576 4252 1584
rect 4074 1500 4194 1506
rect 3857 752 3915 753
rect 4007 752 4045 1458
rect 4074 1392 4080 1500
rect 4188 1392 4194 1500
rect 4074 1386 4194 1392
rect 3857 664 4045 752
rect 4136 717 4197 755
rect 3857 658 4126 664
rect 3857 514 3942 658
rect 4110 514 4126 658
rect 3857 508 4126 514
rect 3857 420 4045 508
rect 4159 461 4197 717
rect 4139 423 4197 461
rect 4233 714 4292 752
rect 4233 465 4271 714
rect 4383 664 4421 1585
rect 4562 1576 4628 1588
rect 4656 1551 4694 1590
rect 4862 1551 4874 1603
rect 4938 1588 4950 1630
rect 4992 1588 5004 1630
rect 5314 1630 5380 1653
rect 4938 1576 5004 1588
rect 5058 1603 5250 1610
rect 4656 1548 4874 1551
rect 4632 1544 4874 1548
rect 5058 1551 5070 1603
rect 5238 1551 5250 1603
rect 5314 1588 5326 1630
rect 5368 1588 5380 1630
rect 5314 1576 5380 1588
rect 5690 1630 5756 1653
rect 5690 1588 5702 1630
rect 5744 1588 5756 1630
rect 5058 1544 5250 1551
rect 4452 1500 4572 1506
rect 4452 1392 4458 1500
rect 4566 1392 4572 1500
rect 4632 1458 4797 1544
rect 4452 1386 4572 1392
rect 4759 754 4797 1458
rect 4886 1498 5048 1504
rect 4886 1402 4892 1498
rect 5042 1402 5048 1498
rect 4886 1396 5048 1402
rect 4610 753 4797 754
rect 4512 714 4573 752
rect 4302 658 4502 664
rect 4302 514 4318 658
rect 4486 514 4502 658
rect 4302 508 4502 514
rect 4233 427 4291 465
rect 3857 419 3916 420
rect 3204 54 3274 60
rect 3370 -378 3608 54
rect 3731 -360 3743 -156
rect 3836 -234 3958 -224
rect 3836 -334 3846 -234
rect 3946 -286 3958 -234
rect 4007 -286 4045 420
rect 4212 -234 4334 -224
rect 3946 -334 4046 -286
rect 3836 -344 4046 -334
rect 4212 -334 4222 -234
rect 4322 -334 4334 -234
rect 4212 -344 4334 -334
rect 3204 -384 3274 -378
rect 3712 -484 3762 -360
rect 3880 -412 4046 -344
rect 4007 -415 4045 -412
rect 4383 -415 4421 508
rect 4535 459 4573 714
rect 4515 421 4573 459
rect 4609 664 4797 753
rect 4888 715 5044 752
rect 4888 714 5021 715
rect 4609 657 4874 664
rect 4609 515 4694 657
rect 4862 515 4874 657
rect 4609 508 4874 515
rect 4609 422 4798 508
rect 4909 459 5021 714
rect 5135 664 5173 1544
rect 5264 714 5327 752
rect 5058 657 5250 664
rect 5058 515 5070 657
rect 5238 515 5250 657
rect 5058 508 5250 515
rect 4909 457 5045 459
rect 4609 421 4797 422
rect 4610 420 4797 421
rect 4607 -286 4668 -284
rect 4759 -286 4797 420
rect 4885 421 5045 457
rect 4885 419 5020 421
rect 4910 418 5020 419
rect 4607 -374 4798 -286
rect 4888 -322 5041 -284
rect 5135 -374 5173 508
rect 5289 459 5327 714
rect 5265 421 5327 459
rect 5361 715 5420 753
rect 5361 459 5399 715
rect 5511 662 5549 1587
rect 5690 1576 5756 1588
rect 5640 1456 5795 1494
rect 5731 751 5796 752
rect 5637 744 5796 751
rect 5637 713 5668 744
rect 5436 657 5624 662
rect 5436 515 5446 657
rect 5614 515 5624 657
rect 5436 510 5624 515
rect 5361 421 5421 459
rect 5204 -218 5326 -210
rect 5204 -322 5214 -218
rect 5316 -322 5326 -218
rect 5204 -330 5326 -322
rect 4607 -420 5250 -374
rect 3498 -530 4502 -484
rect 3498 -608 3670 -530
rect 3204 -656 3258 -640
rect 3204 -698 3210 -656
rect 3252 -658 3258 -656
rect 3252 -696 3449 -658
rect 3252 -698 3258 -696
rect 3204 -716 3258 -698
rect 3212 -723 3250 -716
rect 3204 -913 3258 -897
rect 3204 -955 3210 -913
rect 3252 -915 3258 -913
rect 3411 -915 3449 -696
rect 3631 -912 3670 -608
rect 3836 -574 3956 -564
rect 3836 -674 3846 -574
rect 3946 -674 3956 -574
rect 3836 -684 3956 -674
rect 3480 -913 3670 -912
rect 3252 -953 3449 -915
rect 3252 -955 3258 -953
rect 3204 -973 3258 -955
rect 3212 -979 3250 -973
rect 3204 -1170 3258 -1154
rect 3204 -1212 3210 -1170
rect 3252 -1172 3258 -1170
rect 3411 -1172 3449 -953
rect 3252 -1210 3449 -1172
rect 3252 -1212 3258 -1210
rect 3204 -1230 3258 -1212
rect 3212 -1236 3250 -1230
rect 3204 -1428 3258 -1412
rect 3204 -1470 3210 -1428
rect 3252 -1430 3258 -1428
rect 3411 -1430 3449 -1210
rect 3479 -994 3670 -913
rect 3760 -951 3821 -913
rect 3479 -1000 3750 -994
rect 3479 -1142 3566 -1000
rect 3734 -1142 3750 -1000
rect 3479 -1148 3750 -1142
rect 3479 -1226 3670 -1148
rect 3783 -1193 3821 -951
rect 3479 -1228 3540 -1226
rect 3252 -1468 3449 -1430
rect 3252 -1470 3258 -1468
rect 3204 -1488 3258 -1470
rect 3404 -1478 3449 -1468
rect 3404 -1484 3456 -1478
rect 3212 -1494 3250 -1488
rect 3631 -1532 3670 -1226
rect 3761 -1231 3821 -1193
rect 3857 -952 3916 -914
rect 3857 -1193 3895 -952
rect 4007 -994 4045 -530
rect 4212 -574 4332 -564
rect 4212 -674 4222 -574
rect 4322 -674 4332 -574
rect 4212 -684 4332 -674
rect 4136 -952 4197 -914
rect 3926 -1000 4126 -994
rect 3926 -1142 3942 -1000
rect 4110 -1142 4126 -1000
rect 3926 -1148 4126 -1142
rect 3857 -1231 3917 -1193
rect 3404 -1542 3456 -1536
rect 3498 -1612 3670 -1532
rect 3698 -1466 3818 -1460
rect 3698 -1574 3704 -1466
rect 3812 -1574 3818 -1466
rect 3698 -1580 3818 -1574
rect 4007 -1612 4045 -1148
rect 4159 -1193 4197 -952
rect 4137 -1231 4197 -1193
rect 4233 -951 4292 -913
rect 4233 -1191 4271 -951
rect 4383 -994 4421 -530
rect 4607 -573 4645 -420
rect 4607 -611 4667 -573
rect 4512 -952 4571 -914
rect 4302 -1000 4502 -994
rect 4302 -1142 4318 -1000
rect 4486 -1142 4502 -1000
rect 4302 -1148 4502 -1142
rect 4233 -1229 4291 -1191
rect 4074 -1466 4194 -1460
rect 4074 -1574 4080 -1466
rect 4188 -1574 4194 -1466
rect 4074 -1580 4194 -1574
rect 4383 -1612 4421 -1148
rect 4533 -1191 4571 -952
rect 4513 -1229 4571 -1191
rect 4609 -951 4669 -913
rect 4609 -1190 4647 -951
rect 4759 -994 4797 -488
rect 4888 -610 5045 -572
rect 4888 -932 5044 -914
rect 4888 -952 4925 -932
rect 4682 -1000 4874 -994
rect 4682 -1142 4694 -1000
rect 4862 -1142 4874 -1000
rect 4682 -1148 4874 -1142
rect 4609 -1228 4668 -1190
rect 4450 -1466 4570 -1460
rect 4450 -1574 4456 -1466
rect 4564 -1574 4570 -1466
rect 4450 -1580 4570 -1574
rect 3498 -1618 3750 -1612
rect 3498 -1658 3566 -1618
rect 3550 -1670 3566 -1658
rect 3734 -1670 3750 -1618
rect 3550 -1676 3750 -1670
rect 3926 -1618 4126 -1612
rect 3926 -1670 3942 -1618
rect 4110 -1670 4126 -1618
rect 3926 -1676 4126 -1670
rect 4302 -1618 4502 -1612
rect 4302 -1670 4318 -1618
rect 4486 -1670 4502 -1618
rect 4759 -1653 4797 -1148
rect 4909 -1191 4925 -952
rect 4889 -1212 4925 -1191
rect 5005 -952 5044 -932
rect 5005 -1189 5021 -952
rect 5135 -994 5173 -489
rect 5288 -564 5326 -330
rect 5204 -574 5326 -564
rect 5204 -676 5214 -574
rect 5316 -676 5326 -574
rect 5361 -321 5420 -283
rect 5361 -484 5399 -321
rect 5511 -413 5549 510
rect 5661 458 5668 713
rect 5640 428 5668 458
rect 5762 714 5796 744
rect 5762 604 5769 714
rect 5887 657 5925 1583
rect 6016 714 6075 752
rect 5762 566 5771 604
rect 5762 457 5769 566
rect 5762 428 5791 457
rect 5640 420 5791 428
rect 5731 419 5791 420
rect 5640 -322 5795 -284
rect 5887 -415 5925 515
rect 6037 457 6075 714
rect 6017 419 6075 457
rect 5966 -220 6086 -212
rect 5966 -324 5976 -220
rect 6078 -324 6086 -220
rect 5966 -332 6086 -324
rect 5361 -488 5550 -484
rect 5361 -526 5927 -488
rect 5361 -611 5550 -526
rect 5640 -610 5795 -572
rect 5362 -612 5550 -611
rect 5204 -684 5326 -676
rect 5511 -914 5549 -612
rect 5264 -952 5323 -914
rect 5058 -1000 5250 -994
rect 5058 -1142 5070 -1000
rect 5238 -1142 5250 -1000
rect 5058 -1148 5250 -1142
rect 5005 -1212 5043 -1189
rect 4889 -1227 5043 -1212
rect 4889 -1228 5020 -1227
rect 4888 -1570 5043 -1532
rect 5135 -1654 5173 -1148
rect 5285 -1193 5323 -952
rect 5265 -1231 5323 -1193
rect 5359 -992 5549 -914
rect 5640 -952 5796 -914
rect 5359 -1000 5626 -992
rect 5359 -1142 5446 -1000
rect 5614 -1142 5626 -1000
rect 5359 -1148 5626 -1142
rect 5359 -1228 5549 -1148
rect 5663 -1191 5776 -952
rect 5887 -994 5925 -526
rect 6047 -562 6086 -332
rect 5966 -570 6086 -562
rect 5966 -674 5976 -570
rect 6078 -674 6086 -570
rect 5966 -684 6086 -674
rect 6016 -952 6075 -914
rect 5810 -1000 6002 -994
rect 5810 -1142 5822 -1000
rect 5990 -1142 6002 -1000
rect 5810 -1148 6002 -1142
rect 5663 -1193 5795 -1191
rect 5359 -1229 5419 -1228
rect 5382 -1534 5420 -1532
rect 5511 -1534 5549 -1228
rect 5643 -1229 5795 -1193
rect 5643 -1230 5776 -1229
rect 5636 -1460 5800 -1454
rect 5382 -1604 5550 -1534
rect 5636 -1568 5642 -1460
rect 5794 -1568 5800 -1460
rect 5636 -1574 5800 -1568
rect 5887 -1604 5925 -1148
rect 6037 -1189 6075 -952
rect 6017 -1227 6075 -1189
rect 5382 -1610 5620 -1604
rect 5382 -1653 5446 -1610
rect 5440 -1662 5446 -1653
rect 5614 -1662 5620 -1610
rect 5440 -1668 5620 -1662
rect 5816 -1610 5996 -1604
rect 5816 -1662 5822 -1610
rect 5990 -1662 5996 -1610
rect 5816 -1668 5996 -1662
rect 4302 -1676 4502 -1670
<< via1 >>
rect 4193 1630 4245 1636
rect 4193 1588 4198 1630
rect 4198 1588 4240 1630
rect 4240 1588 4245 1630
rect 4193 1584 4245 1588
rect 4080 1392 4188 1500
rect 3942 514 4110 658
rect 4694 1551 4862 1603
rect 5070 1551 5238 1603
rect 4458 1392 4566 1500
rect 4892 1402 5042 1498
rect 4318 514 4486 658
rect 3204 -378 3274 54
rect 3846 -334 3946 -234
rect 4222 -334 4322 -234
rect 4694 515 4862 657
rect 5070 515 5238 657
rect 5446 515 5614 657
rect 5214 -322 5316 -218
rect 3846 -674 3946 -574
rect 3566 -1142 3734 -1000
rect 3404 -1536 3456 -1484
rect 4222 -674 4322 -574
rect 3942 -1142 4110 -1000
rect 3704 -1574 3812 -1466
rect 4318 -1142 4486 -1000
rect 4080 -1574 4188 -1466
rect 4694 -1142 4862 -1000
rect 4456 -1574 4564 -1466
rect 3566 -1670 3734 -1618
rect 3942 -1670 4110 -1618
rect 4318 -1670 4486 -1618
rect 4925 -1212 5005 -932
rect 5214 -676 5316 -574
rect 5668 428 5762 744
rect 5822 515 5990 657
rect 5976 -324 6078 -220
rect 5070 -1142 5238 -1000
rect 5446 -1142 5614 -1000
rect 5976 -674 6078 -570
rect 5822 -1142 5990 -1000
rect 5642 -1568 5794 -1460
rect 5446 -1662 5614 -1610
rect 5822 -1662 5990 -1610
<< metal2 >>
rect 4187 1584 4193 1636
rect 4245 1584 4251 1636
rect 4682 1603 5250 1610
rect 4194 1506 4244 1584
rect 4682 1551 4694 1603
rect 4862 1551 5070 1603
rect 5238 1551 5250 1603
rect 4682 1546 5250 1551
rect 4074 1500 4274 1506
rect 4074 1474 4080 1500
rect 4188 1496 4274 1500
rect 3214 1426 4080 1474
rect 3214 60 3262 1426
rect 4074 1392 4080 1426
rect 4264 1474 4274 1496
rect 4452 1500 4652 1506
rect 4452 1474 4458 1500
rect 4566 1496 4652 1500
rect 4264 1426 4458 1474
rect 4074 1316 4084 1392
rect 4264 1316 4274 1426
rect 4074 1306 4274 1316
rect 4452 1392 4458 1426
rect 4642 1474 4652 1496
rect 4864 1498 5064 1504
rect 4864 1494 4892 1498
rect 5042 1494 5064 1498
rect 4864 1474 4874 1494
rect 4642 1426 4874 1474
rect 4452 1316 4462 1392
rect 4642 1316 4652 1426
rect 4452 1306 4652 1316
rect 4864 1314 4874 1426
rect 5054 1314 5064 1494
rect 4864 1304 5064 1314
rect 4558 806 5739 854
rect 3926 658 4126 664
rect 3926 514 3942 658
rect 4110 611 4126 658
rect 4302 658 4502 664
rect 4302 611 4318 658
rect 4110 561 4318 611
rect 4110 514 4126 561
rect 3926 508 4126 514
rect 4302 514 4318 561
rect 4486 514 4502 658
rect 4302 508 4502 514
rect 3204 54 3274 60
rect 3836 -234 3958 -224
rect 3836 -334 3846 -234
rect 3946 -334 3958 -234
rect 3836 -344 3958 -334
rect 4212 -234 4334 -224
rect 4212 -334 4222 -234
rect 4322 -260 4334 -234
rect 4558 -260 4606 806
rect 5691 750 5739 806
rect 5662 744 5768 750
rect 4682 657 4874 664
rect 4682 515 4694 657
rect 4862 611 4874 657
rect 5058 657 5250 664
rect 5058 611 5070 657
rect 4862 561 5070 611
rect 4862 515 4874 561
rect 4682 508 4874 515
rect 5058 515 5070 561
rect 5238 515 5250 657
rect 5058 508 5250 515
rect 5436 657 5624 662
rect 5436 515 5446 657
rect 5614 515 5624 657
rect 5436 510 5624 515
rect 5506 178 5554 510
rect 5662 428 5668 744
rect 5762 428 5768 744
rect 5810 657 6002 662
rect 5810 515 5822 657
rect 5990 515 6002 657
rect 5810 510 6002 515
rect 5662 422 5768 428
rect 4322 -308 4606 -260
rect 4752 130 5554 178
rect 4322 -334 4334 -308
rect 4212 -344 4334 -334
rect 3204 -384 3274 -378
rect 3214 -448 3264 -384
rect 3204 -458 3404 -448
rect 3204 -638 3214 -458
rect 3394 -638 3404 -458
rect 3871 -564 3921 -344
rect 4752 -430 4800 130
rect 5882 -32 5930 510
rect 4116 -478 4800 -430
rect 3204 -648 3404 -638
rect 3836 -574 3956 -564
rect 3836 -674 3846 -574
rect 3946 -674 3956 -574
rect 3836 -684 3956 -674
rect 3204 -760 3404 -706
rect 4116 -760 4164 -478
rect 4212 -574 4332 -564
rect 4212 -674 4222 -574
rect 4322 -598 4332 -574
rect 4322 -646 4614 -598
rect 4322 -674 4332 -646
rect 4212 -684 4332 -674
rect 3204 -808 4164 -760
rect 3204 -906 3404 -808
rect 3204 -1070 3404 -962
rect 3550 -1000 3750 -994
rect 3204 -1118 3492 -1070
rect 3204 -1162 3404 -1118
rect 3204 -1349 3404 -1222
rect 3444 -1262 3492 -1118
rect 3550 -1142 3566 -1000
rect 3734 -1046 3750 -1000
rect 3926 -1000 4126 -994
rect 3926 -1046 3942 -1000
rect 3734 -1096 3942 -1046
rect 3734 -1142 3750 -1096
rect 3550 -1148 3750 -1142
rect 3926 -1142 3942 -1096
rect 4110 -1046 4126 -1000
rect 4302 -1000 4502 -994
rect 4302 -1046 4318 -1000
rect 4110 -1096 4318 -1046
rect 4110 -1142 4126 -1096
rect 3926 -1148 4126 -1142
rect 4302 -1142 4318 -1096
rect 4486 -1142 4502 -1000
rect 4302 -1148 4502 -1142
rect 4566 -1178 4614 -646
rect 4752 -994 4800 -478
rect 5128 -80 5930 -32
rect 4909 -932 5021 -914
rect 4682 -1000 4874 -994
rect 4682 -1142 4694 -1000
rect 4862 -1142 4874 -1000
rect 4682 -1148 4874 -1142
rect 4909 -1178 4925 -932
rect 4566 -1212 4925 -1178
rect 5005 -1212 5021 -932
rect 5128 -994 5176 -80
rect 5204 -218 5326 -210
rect 5204 -322 5214 -218
rect 5316 -322 5326 -218
rect 5204 -330 5326 -322
rect 5932 -220 6132 -130
rect 5932 -324 5976 -220
rect 6078 -324 6132 -220
rect 5932 -330 6132 -324
rect 5240 -427 5290 -330
rect 6002 -427 6052 -330
rect 5240 -477 6052 -427
rect 5240 -564 5290 -477
rect 6002 -562 6052 -477
rect 5204 -574 5326 -564
rect 5204 -676 5214 -574
rect 5316 -676 5326 -574
rect 5204 -684 5326 -676
rect 5966 -570 6086 -562
rect 5966 -674 5976 -570
rect 6078 -674 6086 -570
rect 5966 -684 6086 -674
rect 5240 -865 5290 -684
rect 5240 -915 5337 -865
rect 5058 -1000 5250 -994
rect 5058 -1142 5070 -1000
rect 5238 -1142 5250 -1000
rect 5058 -1148 5250 -1142
rect 4566 -1226 5021 -1212
rect 5130 -1262 5178 -1148
rect 3444 -1310 5178 -1262
rect 5287 -1349 5337 -915
rect 5432 -1000 5626 -992
rect 5432 -1142 5446 -1000
rect 5614 -1046 5626 -1000
rect 5810 -1000 6002 -994
rect 5810 -1046 5822 -1000
rect 5614 -1096 5822 -1046
rect 5614 -1142 5626 -1096
rect 5432 -1148 5626 -1142
rect 5810 -1142 5822 -1096
rect 5990 -1142 6002 -1000
rect 5810 -1148 6002 -1142
rect 3204 -1399 5337 -1349
rect 3204 -1422 3404 -1399
rect 3624 -1440 3888 -1430
rect 3204 -1486 3404 -1476
rect 3204 -1666 3214 -1486
rect 3394 -1536 3404 -1486
rect 3456 -1490 3462 -1484
rect 3624 -1490 3634 -1440
rect 3456 -1536 3634 -1490
rect 3394 -1538 3634 -1536
rect 3394 -1666 3404 -1538
rect 3624 -1572 3634 -1538
rect 3878 -1490 3888 -1440
rect 4000 -1438 4264 -1428
rect 4000 -1490 4010 -1438
rect 3878 -1538 4010 -1490
rect 3878 -1572 3888 -1538
rect 3624 -1574 3704 -1572
rect 3812 -1574 3888 -1572
rect 3624 -1582 3888 -1574
rect 4000 -1570 4010 -1538
rect 4254 -1490 4264 -1438
rect 4376 -1438 4640 -1428
rect 4376 -1490 4386 -1438
rect 4254 -1538 4386 -1490
rect 4254 -1570 4264 -1538
rect 4000 -1574 4080 -1570
rect 4188 -1574 4264 -1570
rect 4000 -1580 4264 -1574
rect 4376 -1570 4386 -1538
rect 4630 -1490 4640 -1438
rect 5584 -1434 5848 -1424
rect 5584 -1490 5594 -1434
rect 4630 -1538 5594 -1490
rect 4630 -1570 4640 -1538
rect 4376 -1574 4456 -1570
rect 4564 -1574 4640 -1570
rect 4376 -1580 4640 -1574
rect 5584 -1566 5594 -1538
rect 5838 -1566 5848 -1434
rect 5584 -1568 5642 -1566
rect 5794 -1568 5848 -1566
rect 5584 -1576 5848 -1568
rect 5434 -1610 5630 -1604
rect 5806 -1610 6004 -1604
rect 3204 -1676 3404 -1666
rect 3550 -1618 3750 -1612
rect 3550 -1670 3566 -1618
rect 3734 -1619 3750 -1618
rect 3926 -1618 4126 -1612
rect 3926 -1619 3942 -1618
rect 3734 -1669 3942 -1619
rect 3734 -1670 3750 -1669
rect 3550 -1676 3750 -1670
rect 3926 -1670 3942 -1669
rect 4110 -1619 4126 -1618
rect 4302 -1618 4502 -1612
rect 4302 -1619 4318 -1618
rect 4110 -1669 4318 -1619
rect 4110 -1670 4126 -1669
rect 3926 -1676 4126 -1670
rect 4302 -1670 4318 -1669
rect 4486 -1670 4502 -1618
rect 5434 -1662 5446 -1610
rect 5614 -1660 5822 -1610
rect 5614 -1662 5630 -1660
rect 5434 -1668 5630 -1662
rect 5806 -1662 5822 -1660
rect 5990 -1662 6004 -1610
rect 5806 -1668 6004 -1662
rect 4302 -1676 4502 -1670
<< via2 >>
rect 4084 1392 4188 1496
rect 4188 1392 4264 1496
rect 4084 1316 4264 1392
rect 4462 1392 4566 1496
rect 4566 1392 4642 1496
rect 4462 1316 4642 1392
rect 4874 1402 4892 1494
rect 4892 1402 5042 1494
rect 5042 1402 5054 1494
rect 4874 1314 5054 1402
rect 3214 -638 3394 -458
rect 3214 -1666 3394 -1486
rect 3634 -1466 3878 -1440
rect 3634 -1572 3704 -1466
rect 3704 -1572 3812 -1466
rect 3812 -1572 3878 -1466
rect 4010 -1466 4254 -1438
rect 4010 -1570 4080 -1466
rect 4080 -1570 4188 -1466
rect 4188 -1570 4254 -1466
rect 4386 -1466 4630 -1438
rect 4386 -1570 4456 -1466
rect 4456 -1570 4564 -1466
rect 4564 -1570 4630 -1466
rect 5594 -1460 5838 -1434
rect 5594 -1566 5642 -1460
rect 5642 -1566 5794 -1460
rect 5794 -1566 5838 -1460
<< metal3 >>
rect 4074 1496 4274 1506
rect 4074 1316 4084 1496
rect 4264 1316 4274 1496
rect 4074 688 4274 1316
rect 4452 1496 4652 1506
rect 4452 1316 4462 1496
rect 4642 1316 4652 1496
rect 4452 688 4652 1316
rect 4864 1494 5064 1504
rect 4864 1314 4874 1494
rect 5054 1314 5064 1494
rect 4864 688 5064 1314
rect 3856 488 6074 688
rect 3204 -458 3404 -448
rect 3204 -638 3214 -458
rect 3394 -638 3404 -458
rect 3204 -648 3404 -638
rect 3480 -1162 6074 -962
rect 3656 -1430 3856 -1162
rect 4032 -1428 4232 -1162
rect 4408 -1428 4608 -1162
rect 5616 -1424 5816 -1162
rect 3624 -1440 3888 -1430
rect 3204 -1486 3404 -1476
rect 3204 -1666 3214 -1486
rect 3394 -1666 3404 -1486
rect 3624 -1572 3634 -1440
rect 3878 -1572 3888 -1440
rect 3624 -1582 3888 -1572
rect 4000 -1438 4264 -1428
rect 4000 -1570 4010 -1438
rect 4254 -1570 4264 -1438
rect 4000 -1580 4264 -1570
rect 4376 -1438 4640 -1428
rect 4376 -1570 4386 -1438
rect 4630 -1570 4640 -1438
rect 4376 -1580 4640 -1570
rect 5584 -1434 5848 -1424
rect 5584 -1566 5594 -1434
rect 5838 -1566 5848 -1434
rect 5584 -1576 5848 -1566
rect 3656 -1606 3856 -1582
rect 4032 -1604 4232 -1580
rect 4408 -1604 4608 -1580
rect 5616 -1600 5816 -1576
rect 3204 -1676 3404 -1666
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_0 cells
timestamp 1713334679
transform 1 0 5906 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_1
timestamp 1713334679
transform 1 0 3650 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_2
timestamp 1713334679
transform 1 0 4026 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_3
timestamp 1713334679
transform 1 0 4402 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_4
timestamp 1713334679
transform 1 0 4778 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_5
timestamp 1713334679
transform 1 0 5154 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__nfet_g5v0d10v5_H94GUP  sky130_fd_pr__nfet_g5v0d10v5_H94GUP_6
timestamp 1713334679
transform 1 0 5530 0 1 -1071
box -158 -597 158 597
use sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ  sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ_0 cells
timestamp 1713334679
transform 1 0 4778 0 1 586
box -224 -1018 224 1018
use sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ  sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ_1
timestamp 1713334679
transform 1 0 4026 0 1 586
box -224 -1018 224 1018
use sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ  sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ_2
timestamp 1713334679
transform 1 0 4402 0 1 586
box -224 -1018 224 1018
use sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ  sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ_3
timestamp 1713334679
transform 1 0 5530 0 1 586
box -224 -1018 224 1018
use sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ  sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ_4
timestamp 1713334679
transform 1 0 5154 0 1 586
box -224 -1018 224 1018
use sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ  sky130_fd_pr__pfet_g5v0d10v5_EFU7LQ_5
timestamp 1713334679
transform 1 0 5906 0 1 586
box -224 -1018 224 1018
use sky130_fd_pr__res_xhigh_po_0p35_MDZYBC  sky130_fd_pr__res_xhigh_po_0p35_MDZYBC_0 cells
timestamp 1713341356
transform 1 0 3488 0 -1 663
box -284 -1041 284 1041
<< labels >>
flabel metal2 5932 -330 6132 -130 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal3 3204 -648 3404 -448 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal2 3204 -906 3404 -706 0 FreeSans 256 0 0 0 P
port 2 nsew
flabel metal2 3204 -1162 3404 -962 0 FreeSans 256 0 0 0 N
port 3 nsew
flabel metal2 3204 -1422 3404 -1222 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal3 4864 1304 5064 1504 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 3624 -1582 3888 -1430 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal3 4000 -1580 4264 -1428 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal3 4376 -1580 4640 -1428 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal3 5584 -1576 5848 -1424 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal3 3856 488 6074 688 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 3480 -1162 6074 -962 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal3 4452 1306 4652 1506 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 4074 1306 4274 1506 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 3204 -1676 3404 -1476 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
