magic
tech sky130A
magscale 1 2
timestamp 1762787048
<< metal1 >>
rect 2820 42702 3220 42708
rect 3220 42302 4732 42702
rect 2820 42296 3220 42302
rect 25016 41454 25348 41460
rect 23792 41122 25016 41454
rect 25016 41116 25348 41122
rect 23422 39504 23428 39564
rect 23488 39504 23494 39564
rect 23428 38890 23488 39504
rect 3146 35280 3546 35286
rect 3546 34880 4634 35280
rect 3146 34874 3546 34880
<< via1 >>
rect 2820 42302 3220 42702
rect 25016 41122 25348 41454
rect 23428 39504 23488 39564
rect 3146 34880 3546 35280
<< metal2 >>
rect 1949 42702 2339 42706
rect 1944 42697 2820 42702
rect 1944 42307 1949 42697
rect 2339 42307 2820 42697
rect 1944 42302 2820 42307
rect 3220 42302 3226 42702
rect 1949 42298 2339 42302
rect 25010 41122 25016 41454
rect 25348 41122 25354 41454
rect 23428 39694 23488 39696
rect 23421 39638 23430 39694
rect 23486 39638 23495 39694
rect 23428 39564 23488 39638
rect 23428 39498 23488 39504
rect 2631 35280 3021 35284
rect 2626 35275 3146 35280
rect 2626 34885 2631 35275
rect 3021 34885 3146 35275
rect 2626 34880 3146 34885
rect 3546 34880 3552 35280
rect 2631 34876 3021 34880
rect 25016 3228 25348 41122
rect 26092 3964 26626 3973
rect 26092 3318 26626 3430
rect 25074 3058 25291 3228
rect 26076 3130 27084 3318
rect 25074 2874 27100 3058
rect 25074 2858 25291 2874
rect 26136 2608 27106 2808
rect 26136 2558 26336 2608
rect 26136 2358 27100 2558
rect 26186 1197 26366 2358
rect 26666 1674 27126 2264
rect 26611 1670 27126 1674
rect 26606 1665 27232 1670
rect 26606 1275 26611 1665
rect 27001 1275 27232 1665
rect 26606 1270 27232 1275
rect 26611 1266 27001 1270
rect 26182 1027 26191 1197
rect 26361 1027 26370 1197
rect 26186 1022 26366 1027
<< via2 >>
rect 1949 42307 2339 42697
rect 23430 39638 23486 39694
rect 2631 34885 3021 35275
rect 26092 3430 26626 3964
rect 26611 1275 27001 1665
rect 26191 1027 26361 1197
<< metal3 >>
rect 190 42702 606 42712
rect 190 42701 2344 42702
rect 190 42303 201 42701
rect 599 42697 2344 42701
rect 599 42307 1949 42697
rect 2339 42307 2344 42697
rect 599 42303 2344 42307
rect 190 42302 2344 42303
rect 190 42294 606 42302
rect 23426 39910 23490 39916
rect 23426 39840 23490 39846
rect 23428 39699 23488 39840
rect 23425 39694 23491 39699
rect 23425 39638 23430 39694
rect 23486 39638 23491 39694
rect 23425 39633 23491 39638
rect 1833 35280 2231 35285
rect 1832 35279 3026 35280
rect 1832 34881 1833 35279
rect 2231 35275 3026 35279
rect 2231 34885 2631 35275
rect 3021 34885 3026 35275
rect 2231 34881 3026 34885
rect 1832 34880 3026 34881
rect 1833 34875 2231 34880
rect 23887 4173 26626 4707
rect 3664 2562 4092 2582
rect 214 2526 4092 2562
rect 214 2216 230 2526
rect 578 2216 4092 2526
rect 214 2174 4092 2216
rect 3664 1138 4092 2174
rect 23940 1138 24368 4173
rect 26092 3969 26626 4173
rect 26087 3964 26631 3969
rect 26087 3430 26092 3964
rect 26626 3430 26631 3964
rect 26087 3425 26631 3430
rect 24891 1670 25289 1675
rect 24890 1669 27006 1670
rect 24890 1271 24891 1669
rect 25289 1665 27006 1669
rect 25289 1275 26611 1665
rect 27001 1275 27006 1665
rect 25289 1271 27006 1275
rect 24890 1270 27006 1271
rect 24891 1265 25289 1270
rect 3664 710 24368 1138
rect 26186 1197 26366 1202
rect 26186 1027 26191 1197
rect 26361 1027 26366 1197
rect 26186 961 26366 1027
rect 26181 783 26187 961
rect 26365 783 26371 961
rect 26186 782 26366 783
<< via3 >>
rect 201 42303 599 42701
rect 23426 39846 23490 39910
rect 1833 34881 2231 35279
rect 230 2216 578 2526
rect 24891 1271 25289 1669
rect 26187 783 26365 961
<< metal4 >>
rect 200 42701 600 44152
rect 200 42303 201 42701
rect 599 42303 600 42701
rect 200 2526 600 42303
rect 200 2216 230 2526
rect 578 2216 600 2526
rect 200 1000 600 2216
rect 800 44002 1200 44152
rect 6134 44002 6194 45152
rect 6686 44002 6746 45152
rect 7238 44002 7298 45152
rect 7790 44002 7850 45152
rect 8342 44002 8402 45152
rect 8894 44002 8954 45152
rect 9446 44002 9506 45152
rect 9998 44002 10058 45152
rect 10550 44002 10610 45152
rect 11102 44002 11162 45152
rect 11654 44002 11714 45152
rect 12206 44002 12266 45152
rect 12758 44002 12818 45152
rect 13310 44002 13370 45152
rect 13862 44002 13922 45152
rect 14414 44002 14474 45152
rect 14966 44002 15026 45152
rect 15518 44002 15578 45152
rect 16070 44002 16130 45152
rect 16622 44002 16682 45152
rect 17174 44002 17234 45152
rect 17726 44002 17786 45152
rect 18278 44002 18338 45152
rect 18830 44286 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 18830 44226 23488 44286
rect 800 43602 18486 44002
rect 800 35280 1200 43602
rect 23428 39911 23488 44226
rect 23425 39910 23491 39911
rect 23425 39846 23426 39910
rect 23490 39846 23491 39910
rect 23425 39845 23491 39846
rect 800 35279 2232 35280
rect 800 34881 1833 35279
rect 2231 34881 2232 35279
rect 800 34880 2232 34881
rect 800 1670 1200 34880
rect 800 1669 25290 1670
rect 800 1271 24891 1669
rect 25289 1271 25290 1669
rect 800 1270 25290 1271
rect 800 1000 1200 1270
rect 26186 961 30542 962
rect 26186 783 26187 961
rect 26365 783 30542 961
rect 26186 782 30542 783
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 782
use osc  osc_0
timestamp 1762786006
transform 1 0 -308 0 1 29588
box 3800 -27612 24528 13400
use vfollower  vfollower_0
timestamp 1713341356
transform 1 0 26538 0 1 3292
box 368 -1198 3296 2198
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
